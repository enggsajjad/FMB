library verilog;
use verilog.vl_types.all;
entity tf_top_tx is
end tf_top_tx;
