module test_uart(din_byte,dout_byte);

input [7:0] din_byte;
output [7:0] dout_byte;

assign dout_byte = din_byte;

endmodule
