library verilog;
use verilog.vl_types.all;
entity test_uar_tf is
end test_uar_tf;
